library verilog;
use verilog.vl_types.all;
entity DisplayVal_vlg_vec_tst is
end DisplayVal_vlg_vec_tst;
