library verilog;
use verilog.vl_types.all;
entity procULA_vlg_vec_tst is
end procULA_vlg_vec_tst;
